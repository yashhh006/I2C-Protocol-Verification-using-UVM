`include "i2cSlaveTop.v"
