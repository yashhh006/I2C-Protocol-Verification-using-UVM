`include "top.sv"
