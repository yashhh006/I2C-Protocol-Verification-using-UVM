`ifndef I2C_SQR_SVH
`define I2C_SQR_SVH


typedef uvm_sequencer #(i2c_tx)i2c_sqr;

`endif